`timescale 1 ns / 1 ns

module RXx
          (TB_Encoded_0,
           TB_Encoded_1,
           TB_Encoded_2,
           TB_Encoded_3,
           TB_Encoded_4,
           TB_Encoded_5,
           TB_Encoded_6,
           TB_Encoded_7,
           TB_Encoded_8,
           TB_Encoded_9,
           TB_Encoded_10,
           TB_Encoded_11,
           TB_Encoded_12,
           TB_Encoded_13,
           TB_Encoded_14,
           TB_Encoded_15,
           TB_Encoded_16,
           TB_Encoded_17,
           TB_Encoded_18,
           TB_Encoded_19,
           TB_Encoded_20,
           TB_Encoded_21,
           TB_Encoded_22,
           TB_Encoded_23,
           TB_Encoded_24,
           TB_Encoded_25,
           TB_Encoded_26,
           TB_Encoded_27,
           TB_Encoded_28,
           TB_Encoded_29,
           TB_Encoded_30,
           TB_Encoded_31,
           TB_Encoded_32,
           TB_Encoded_33,
           TB_Encoded_34,
           TB_Encoded_35,
           TB_Encoded_36,
           TB_Encoded_37,
           TB_Encoded_38,
           TB_Encoded_39,
           TB_Encoded_40,
           TB_Encoded_41,
           TB_Encoded_42,
           TB_Encoded_43,
           TB_Encoded_44,
           TB_Encoded_45,
           TB_Encoded_46,
           TB_Encoded_47,
           Lower_zk1_0,
           Lower_zk1_1,
           Lower_zk1_2,
           Lower_zk1_3,
           Lower_zk1_4,
           Lower_zk1_5,
           Lower_zk1_6,
           Lower_zk1_7,
           Lower_zk1_8,
           Lower_zk1_9,
           Lower_zk1_10,
           Lower_zk1_11,
           Lower_zk1_12,
           Lower_zk1_13,
           Lower_zk1_14,
           Lower_zk1_15,
           Lower_zk1_16,
           Lower_zk1_17,
           Lower_zk1_18,
           Lower_zk1_19,
           Lower_zk1_20,
           Lower_zk1_21,
           Lower_zk1_22,
           Lower_zk1_23,
           Lower_zk1_24,
           Lower_zk1_25,
           Lower_zk1_26,
           Lower_zk1_27,
           Lower_zk1_28,
           Lower_zk1_29,
           Lower_zk1_30,
           Lower_zk1_31,
           Lower_zk1_32,
           Lower_zk1_33,
           Lower_zk1_34,
           Lower_zk1_35,
           Lower_zk1_36,
           Lower_zk1_37,
           Lower_zk1_38,
           Lower_zk1_39,
           Lower_zk1_40,
           Lower_zk1_41,
           Lower_zk1_42,
           Lower_zk1_43,
           Lower_zk1_44,
           Lower_zk1_45,
           Lower_zk1_46,
           Lower_zk1_47,
           Upper_zk_0,
           Upper_zk_1,
           Upper_zk_2,
           Upper_zk_3,
           Upper_zk_4,
           Upper_zk_5,
           Upper_zk_6,
           Upper_zk_7,
           Upper_zk_8,
           Upper_zk_9,
           Upper_zk_10,
           Upper_zk_11,
           Upper_zk_12,
           Upper_zk_13,
           Upper_zk_14,
           Upper_zk_15,
           Upper_zk_16,
           Upper_zk_17,
           Upper_zk_18,
           Upper_zk_19,
           Upper_zk_20,
           Upper_zk_21,
           Upper_zk_22,
           Upper_zk_23,
           Upper_zk_24,
           Upper_zk_25,
           Upper_zk_26,
           Upper_zk_27,
           Upper_zk_28,
           Upper_zk_29,
           Upper_zk_30,
           Upper_zk_31,
           Upper_zk_32,
           Upper_zk_33,
           Upper_zk_34,
           Upper_zk_35,
           Upper_zk_36,
           Upper_zk_37,
           Upper_zk_38,
           Upper_zk_39,
           Upper_zk_40,
           Upper_zk_41,
           Upper_zk_42,
           Upper_zk_43,
           Upper_zk_44,
           Upper_zk_45,
           Upper_zk_46,
           Upper_zk_47,
           Final_Decoded_0,
           Final_Decoded_1,
           Final_Decoded_2,
           Final_Decoded_3,
           Final_Decoded_4,
           Final_Decoded_5,
           Final_Decoded_6,
           Final_Decoded_7,
           Final_Decoded_8,
           Final_Decoded_9,
           Final_Decoded_10,
           Final_Decoded_11,
           Final_Decoded_12,
           Final_Decoded_13,
           Final_Decoded_14,
           Final_Decoded_15,
           Final_Decoded_16,
           Final_Decoded_17,
           Final_Decoded_18,
           Final_Decoded_19,
           Final_Decoded_20,
           Final_Decoded_21,
           Final_Decoded_22,
           Final_Decoded_23,
           Final_Decoded_24,
           Final_Decoded_25,
           Final_Decoded_26,
           Final_Decoded_27,
           Final_Decoded_28,
           Final_Decoded_29,
           Final_Decoded_30,
           Final_Decoded_31,
           Final_Decoded_32,
           Final_Decoded_33,
           Final_Decoded_34,
           Final_Decoded_35,
           Final_Decoded_36,
           Final_Decoded_37,
           Final_Decoded_38,
           Final_Decoded_39);


  input   TB_Encoded_0;  // ufix1
  input   TB_Encoded_1;  // ufix1
  input   TB_Encoded_2;  // ufix1
  input   TB_Encoded_3;  // ufix1
  input   TB_Encoded_4;  // ufix1
  input   TB_Encoded_5;  // ufix1
  input   TB_Encoded_6;  // ufix1
  input   TB_Encoded_7;  // ufix1
  input   TB_Encoded_8;  // ufix1
  input   TB_Encoded_9;  // ufix1
  input   TB_Encoded_10;  // ufix1
  input   TB_Encoded_11;  // ufix1
  input   TB_Encoded_12;  // ufix1
  input   TB_Encoded_13;  // ufix1
  input   TB_Encoded_14;  // ufix1
  input   TB_Encoded_15;  // ufix1
  input   TB_Encoded_16;  // ufix1
  input   TB_Encoded_17;  // ufix1
  input   TB_Encoded_18;  // ufix1
  input   TB_Encoded_19;  // ufix1
  input   TB_Encoded_20;  // ufix1
  input   TB_Encoded_21;  // ufix1
  input   TB_Encoded_22;  // ufix1
  input   TB_Encoded_23;  // ufix1
  input   TB_Encoded_24;  // ufix1
  input   TB_Encoded_25;  // ufix1
  input   TB_Encoded_26;  // ufix1
  input   TB_Encoded_27;  // ufix1
  input   TB_Encoded_28;  // ufix1
  input   TB_Encoded_29;  // ufix1
  input   TB_Encoded_30;  // ufix1
  input   TB_Encoded_31;  // ufix1
  input   TB_Encoded_32;  // ufix1
  input   TB_Encoded_33;  // ufix1
  input   TB_Encoded_34;  // ufix1
  input   TB_Encoded_35;  // ufix1
  input   TB_Encoded_36;  // ufix1
  input   TB_Encoded_37;  // ufix1
  input   TB_Encoded_38;  // ufix1
  input   TB_Encoded_39;  // ufix1
  input   TB_Encoded_40;  // ufix1
  input   TB_Encoded_41;  // ufix1
  input   TB_Encoded_42;  // ufix1
  input   TB_Encoded_43;  // ufix1
  input   TB_Encoded_44;  // ufix1
  input   TB_Encoded_45;  // ufix1
  input   TB_Encoded_46;  // ufix1
  input   TB_Encoded_47;  // ufix1
  input   Lower_zk1_0;  // ufix1
  input   Lower_zk1_1;  // ufix1
  input   Lower_zk1_2;  // ufix1
  input   Lower_zk1_3;  // ufix1
  input   Lower_zk1_4;  // ufix1
  input   Lower_zk1_5;  // ufix1
  input   Lower_zk1_6;  // ufix1
  input   Lower_zk1_7;  // ufix1
  input   Lower_zk1_8;  // ufix1
  input   Lower_zk1_9;  // ufix1
  input   Lower_zk1_10;  // ufix1
  input   Lower_zk1_11;  // ufix1
  input   Lower_zk1_12;  // ufix1
  input   Lower_zk1_13;  // ufix1
  input   Lower_zk1_14;  // ufix1
  input   Lower_zk1_15;  // ufix1
  input   Lower_zk1_16;  // ufix1
  input   Lower_zk1_17;  // ufix1
  input   Lower_zk1_18;  // ufix1
  input   Lower_zk1_19;  // ufix1
  input   Lower_zk1_20;  // ufix1
  input   Lower_zk1_21;  // ufix1
  input   Lower_zk1_22;  // ufix1
  input   Lower_zk1_23;  // ufix1
  input   Lower_zk1_24;  // ufix1
  input   Lower_zk1_25;  // ufix1
  input   Lower_zk1_26;  // ufix1
  input   Lower_zk1_27;  // ufix1
  input   Lower_zk1_28;  // ufix1
  input   Lower_zk1_29;  // ufix1
  input   Lower_zk1_30;  // ufix1
  input   Lower_zk1_31;  // ufix1
  input   Lower_zk1_32;  // ufix1
  input   Lower_zk1_33;  // ufix1
  input   Lower_zk1_34;  // ufix1
  input   Lower_zk1_35;  // ufix1
  input   Lower_zk1_36;  // ufix1
  input   Lower_zk1_37;  // ufix1
  input   Lower_zk1_38;  // ufix1
  input   Lower_zk1_39;  // ufix1
  input   Lower_zk1_40;  // ufix1
  input   Lower_zk1_41;  // ufix1
  input   Lower_zk1_42;  // ufix1
  input   Lower_zk1_43;  // ufix1
  input   Lower_zk1_44;  // ufix1
  input   Lower_zk1_45;  // ufix1
  input   Lower_zk1_46;  // ufix1
  input   Lower_zk1_47;  // ufix1
  input   Upper_zk_0;  // ufix1
  input   Upper_zk_1;  // ufix1
  input   Upper_zk_2;  // ufix1
  input   Upper_zk_3;  // ufix1
  input   Upper_zk_4;  // ufix1
  input   Upper_zk_5;  // ufix1
  input   Upper_zk_6;  // ufix1
  input   Upper_zk_7;  // ufix1
  input   Upper_zk_8;  // ufix1
  input   Upper_zk_9;  // ufix1
  input   Upper_zk_10;  // ufix1
  input   Upper_zk_11;  // ufix1
  input   Upper_zk_12;  // ufix1
  input   Upper_zk_13;  // ufix1
  input   Upper_zk_14;  // ufix1
  input   Upper_zk_15;  // ufix1
  input   Upper_zk_16;  // ufix1
  input   Upper_zk_17;  // ufix1
  input   Upper_zk_18;  // ufix1
  input   Upper_zk_19;  // ufix1
  input   Upper_zk_20;  // ufix1
  input   Upper_zk_21;  // ufix1
  input   Upper_zk_22;  // ufix1
  input   Upper_zk_23;  // ufix1
  input   Upper_zk_24;  // ufix1
  input   Upper_zk_25;  // ufix1
  input   Upper_zk_26;  // ufix1
  input   Upper_zk_27;  // ufix1
  input   Upper_zk_28;  // ufix1
  input   Upper_zk_29;  // ufix1
  input   Upper_zk_30;  // ufix1
  input   Upper_zk_31;  // ufix1
  input   Upper_zk_32;  // ufix1
  input   Upper_zk_33;  // ufix1
  input   Upper_zk_34;  // ufix1
  input   Upper_zk_35;  // ufix1
  input   Upper_zk_36;  // ufix1
  input   Upper_zk_37;  // ufix1
  input   Upper_zk_38;  // ufix1
  input   Upper_zk_39;  // ufix1
  input   Upper_zk_40;  // ufix1
  input   Upper_zk_41;  // ufix1
  input   Upper_zk_42;  // ufix1
  input   Upper_zk_43;  // ufix1
  input   Upper_zk_44;  // ufix1
  input   Upper_zk_45;  // ufix1
  input   Upper_zk_46;  // ufix1
  input   Upper_zk_47;  // ufix1
  output  Final_Decoded_0;  // ufix1
  output  Final_Decoded_1;  // ufix1
  output  Final_Decoded_2;  // ufix1
  output  Final_Decoded_3;  // ufix1
  output  Final_Decoded_4;  // ufix1
  output  Final_Decoded_5;  // ufix1
  output  Final_Decoded_6;  // ufix1
  output  Final_Decoded_7;  // ufix1
  output  Final_Decoded_8;  // ufix1
  output  Final_Decoded_9;  // ufix1
  output  Final_Decoded_10;  // ufix1
  output  Final_Decoded_11;  // ufix1
  output  Final_Decoded_12;  // ufix1
  output  Final_Decoded_13;  // ufix1
  output  Final_Decoded_14;  // ufix1
  output  Final_Decoded_15;  // ufix1
  output  Final_Decoded_16;  // ufix1
  output  Final_Decoded_17;  // ufix1
  output  Final_Decoded_18;  // ufix1
  output  Final_Decoded_19;  // ufix1
  output  Final_Decoded_20;  // ufix1
  output  Final_Decoded_21;  // ufix1
  output  Final_Decoded_22;  // ufix1
  output  Final_Decoded_23;  // ufix1
  output  Final_Decoded_24;  // ufix1
  output  Final_Decoded_25;  // ufix1
  output  Final_Decoded_26;  // ufix1
  output  Final_Decoded_27;  // ufix1
  output  Final_Decoded_28;  // ufix1
  output  Final_Decoded_29;  // ufix1
  output  Final_Decoded_30;  // ufix1
  output  Final_Decoded_31;  // ufix1
  output  Final_Decoded_32;  // ufix1
  output  Final_Decoded_33;  // ufix1
  output  Final_Decoded_34;  // ufix1
  output  Final_Decoded_35;  // ufix1
  output  Final_Decoded_36;  // ufix1
  output  Final_Decoded_37;  // ufix1
  output  Final_Decoded_38;  // ufix1
  output  Final_Decoded_39;  // ufix1


  wire [0:47] TB_Encoded;  // ufix1 [48]
  wire [0:47] Lower_zk1;  // ufix1 [48]
  wire [0:47] Upper_zk;  // ufix1 [48]
  reg  [0:39] Final_Decoded;  // ufix1 [40]
  reg signed [1:0] decoder_fun_fixpt_x [0:47];  // sfix2 [48]
  reg  [0:39] decoder_fun_fixpt_Decoded_out;  // ufix1 [40]
  reg [5:0] decoder_fun_fixpt_ii;  // ufix6
  reg signed [2:0] decoder_fun_fixpt_LZ [0:39];  // sfix3 [40]
  reg signed [31:0] decoder_fun_fixpt_ii_0;  // int32
  reg signed [31:0] decoder_fun_fixpt_t_0;  // int32
  reg signed [31:0] decoder_fun_fixpt_t_1;  // int32
  reg signed [4:0] decoder_fun_fixpt_add_cast [0:47];  // sfix5 [48]
  reg signed [4:0] decoder_fun_fixpt_add_temp [0:47];  // sfix5 [48]
  reg signed [31:0] decoder_fun_fixpt_add_temp_0 [0:39];  // int32 [40]
  reg signed [5:0] decoder_fun_fixpt_cast [0:39];  // sfix6 [40]
  reg signed [1:0] decoder_fun_fixpt_t_2 [0:47];  // sfix2 [48]


  assign TB_Encoded[0] = TB_Encoded_0;
  assign TB_Encoded[1] = TB_Encoded_1;
  assign TB_Encoded[2] = TB_Encoded_2;
  assign TB_Encoded[3] = TB_Encoded_3;
  assign TB_Encoded[4] = TB_Encoded_4;
  assign TB_Encoded[5] = TB_Encoded_5;
  assign TB_Encoded[6] = TB_Encoded_6;
  assign TB_Encoded[7] = TB_Encoded_7;
  assign TB_Encoded[8] = TB_Encoded_8;
  assign TB_Encoded[9] = TB_Encoded_9;
  assign TB_Encoded[10] = TB_Encoded_10;
  assign TB_Encoded[11] = TB_Encoded_11;
  assign TB_Encoded[12] = TB_Encoded_12;
  assign TB_Encoded[13] = TB_Encoded_13;
  assign TB_Encoded[14] = TB_Encoded_14;
  assign TB_Encoded[15] = TB_Encoded_15;
  assign TB_Encoded[16] = TB_Encoded_16;
  assign TB_Encoded[17] = TB_Encoded_17;
  assign TB_Encoded[18] = TB_Encoded_18;
  assign TB_Encoded[19] = TB_Encoded_19;
  assign TB_Encoded[20] = TB_Encoded_20;
  assign TB_Encoded[21] = TB_Encoded_21;
  assign TB_Encoded[22] = TB_Encoded_22;
  assign TB_Encoded[23] = TB_Encoded_23;
  assign TB_Encoded[24] = TB_Encoded_24;
  assign TB_Encoded[25] = TB_Encoded_25;
  assign TB_Encoded[26] = TB_Encoded_26;
  assign TB_Encoded[27] = TB_Encoded_27;
  assign TB_Encoded[28] = TB_Encoded_28;
  assign TB_Encoded[29] = TB_Encoded_29;
  assign TB_Encoded[30] = TB_Encoded_30;
  assign TB_Encoded[31] = TB_Encoded_31;
  assign TB_Encoded[32] = TB_Encoded_32;
  assign TB_Encoded[33] = TB_Encoded_33;
  assign TB_Encoded[34] = TB_Encoded_34;
  assign TB_Encoded[35] = TB_Encoded_35;
  assign TB_Encoded[36] = TB_Encoded_36;
  assign TB_Encoded[37] = TB_Encoded_37;
  assign TB_Encoded[38] = TB_Encoded_38;
  assign TB_Encoded[39] = TB_Encoded_39;
  assign TB_Encoded[40] = TB_Encoded_40;
  assign TB_Encoded[41] = TB_Encoded_41;
  assign TB_Encoded[42] = TB_Encoded_42;
  assign TB_Encoded[43] = TB_Encoded_43;
  assign TB_Encoded[44] = TB_Encoded_44;
  assign TB_Encoded[45] = TB_Encoded_45;
  assign TB_Encoded[46] = TB_Encoded_46;
  assign TB_Encoded[47] = TB_Encoded_47;

  assign Lower_zk1[0] = Lower_zk1_0;
  assign Lower_zk1[1] = Lower_zk1_1;
  assign Lower_zk1[2] = Lower_zk1_2;
  assign Lower_zk1[3] = Lower_zk1_3;
  assign Lower_zk1[4] = Lower_zk1_4;
  assign Lower_zk1[5] = Lower_zk1_5;
  assign Lower_zk1[6] = Lower_zk1_6;
  assign Lower_zk1[7] = Lower_zk1_7;
  assign Lower_zk1[8] = Lower_zk1_8;
  assign Lower_zk1[9] = Lower_zk1_9;
  assign Lower_zk1[10] = Lower_zk1_10;
  assign Lower_zk1[11] = Lower_zk1_11;
  assign Lower_zk1[12] = Lower_zk1_12;
  assign Lower_zk1[13] = Lower_zk1_13;
  assign Lower_zk1[14] = Lower_zk1_14;
  assign Lower_zk1[15] = Lower_zk1_15;
  assign Lower_zk1[16] = Lower_zk1_16;
  assign Lower_zk1[17] = Lower_zk1_17;
  assign Lower_zk1[18] = Lower_zk1_18;
  assign Lower_zk1[19] = Lower_zk1_19;
  assign Lower_zk1[20] = Lower_zk1_20;
  assign Lower_zk1[21] = Lower_zk1_21;
  assign Lower_zk1[22] = Lower_zk1_22;
  assign Lower_zk1[23] = Lower_zk1_23;
  assign Lower_zk1[24] = Lower_zk1_24;
  assign Lower_zk1[25] = Lower_zk1_25;
  assign Lower_zk1[26] = Lower_zk1_26;
  assign Lower_zk1[27] = Lower_zk1_27;
  assign Lower_zk1[28] = Lower_zk1_28;
  assign Lower_zk1[29] = Lower_zk1_29;
  assign Lower_zk1[30] = Lower_zk1_30;
  assign Lower_zk1[31] = Lower_zk1_31;
  assign Lower_zk1[32] = Lower_zk1_32;
  assign Lower_zk1[33] = Lower_zk1_33;
  assign Lower_zk1[34] = Lower_zk1_34;
  assign Lower_zk1[35] = Lower_zk1_35;
  assign Lower_zk1[36] = Lower_zk1_36;
  assign Lower_zk1[37] = Lower_zk1_37;
  assign Lower_zk1[38] = Lower_zk1_38;
  assign Lower_zk1[39] = Lower_zk1_39;
  assign Lower_zk1[40] = Lower_zk1_40;
  assign Lower_zk1[41] = Lower_zk1_41;
  assign Lower_zk1[42] = Lower_zk1_42;
  assign Lower_zk1[43] = Lower_zk1_43;
  assign Lower_zk1[44] = Lower_zk1_44;
  assign Lower_zk1[45] = Lower_zk1_45;
  assign Lower_zk1[46] = Lower_zk1_46;
  assign Lower_zk1[47] = Lower_zk1_47;

  assign Upper_zk[0] = Upper_zk_0;
  assign Upper_zk[1] = Upper_zk_1;
  assign Upper_zk[2] = Upper_zk_2;
  assign Upper_zk[3] = Upper_zk_3;
  assign Upper_zk[4] = Upper_zk_4;
  assign Upper_zk[5] = Upper_zk_5;
  assign Upper_zk[6] = Upper_zk_6;
  assign Upper_zk[7] = Upper_zk_7;
  assign Upper_zk[8] = Upper_zk_8;
  assign Upper_zk[9] = Upper_zk_9;
  assign Upper_zk[10] = Upper_zk_10;
  assign Upper_zk[11] = Upper_zk_11;
  assign Upper_zk[12] = Upper_zk_12;
  assign Upper_zk[13] = Upper_zk_13;
  assign Upper_zk[14] = Upper_zk_14;
  assign Upper_zk[15] = Upper_zk_15;
  assign Upper_zk[16] = Upper_zk_16;
  assign Upper_zk[17] = Upper_zk_17;
  assign Upper_zk[18] = Upper_zk_18;
  assign Upper_zk[19] = Upper_zk_19;
  assign Upper_zk[20] = Upper_zk_20;
  assign Upper_zk[21] = Upper_zk_21;
  assign Upper_zk[22] = Upper_zk_22;
  assign Upper_zk[23] = Upper_zk_23;
  assign Upper_zk[24] = Upper_zk_24;
  assign Upper_zk[25] = Upper_zk_25;
  assign Upper_zk[26] = Upper_zk_26;
  assign Upper_zk[27] = Upper_zk_27;
  assign Upper_zk[28] = Upper_zk_28;
  assign Upper_zk[29] = Upper_zk_29;
  assign Upper_zk[30] = Upper_zk_30;
  assign Upper_zk[31] = Upper_zk_31;
  assign Upper_zk[32] = Upper_zk_32;
  assign Upper_zk[33] = Upper_zk_33;
  assign Upper_zk[34] = Upper_zk_34;
  assign Upper_zk[35] = Upper_zk_35;
  assign Upper_zk[36] = Upper_zk_36;
  assign Upper_zk[37] = Upper_zk_37;
  assign Upper_zk[38] = Upper_zk_38;
  assign Upper_zk[39] = Upper_zk_39;
  assign Upper_zk[40] = Upper_zk_40;
  assign Upper_zk[41] = Upper_zk_41;
  assign Upper_zk[42] = Upper_zk_42;
  assign Upper_zk[43] = Upper_zk_43;
  assign Upper_zk[44] = Upper_zk_44;
  assign Upper_zk[45] = Upper_zk_45;
  assign Upper_zk[46] = Upper_zk_46;
  assign Upper_zk[47] = Upper_zk_47;

  always @* begin
    decoder_fun_fixpt_ii = 6'b000000;
    //HDL code generation from MATLAB function: decoder_fun_fixpt
    //+LZ1(1,ii)+LZ2(1,ii);
    //%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%
    //                                                                          %
    //                                                                          %
    //%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%
    //%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%
    //   20(-1)  15(1)  6(-1) 2(1) 1(-1) 4(1)

    for(decoder_fun_fixpt_t_0 = 32'sd0; decoder_fun_fixpt_t_0 <= 32'sd47; decoder_fun_fixpt_t_0 = decoder_fun_fixpt_t_0 + 32'sd1) begin
      if (TB_Encoded[decoder_fun_fixpt_t_0] == 1'b1) begin
        decoder_fun_fixpt_t_2[decoder_fun_fixpt_t_0] = 2'sb10;
      end
      else begin
        decoder_fun_fixpt_t_2[decoder_fun_fixpt_t_0] = 2'sb00;
      end
      decoder_fun_fixpt_add_cast[decoder_fun_fixpt_t_0] = {{3{decoder_fun_fixpt_t_2[decoder_fun_fixpt_t_0][1]}}, decoder_fun_fixpt_t_2[decoder_fun_fixpt_t_0]};
      decoder_fun_fixpt_add_temp[decoder_fun_fixpt_t_0] = decoder_fun_fixpt_add_cast[decoder_fun_fixpt_t_0] + 5'sb00001;
      decoder_fun_fixpt_x[decoder_fun_fixpt_t_0] = decoder_fun_fixpt_add_temp[decoder_fun_fixpt_t_0][1:0];
    end

    //%%%%%%%%%%%%%%%%% Decoder I %%%%%%%%%%%%%%%%%%%%%%%%%%%
    //%%%%%%%%%%%%%%%%% Decoder I END %%%%%%%%%%%%%%%%%%%%%%%%%%%      
    //%%%%%%%%%%%%%%%%% Decoder I alpha forward %%%%%%%%%%%%%%%%%%%%% metr
    //%%%%%%%%%%%%5%%Decoder I beta backward metric%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%
    //%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%     
    //%%%%%interleave the extrensic%%%%%%%%%%%%%%%%%
    //%%%%%%%%%%% Decoder%%% II %%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%
    //%%%%%%%%%%% Decoder%%% II END%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%     
    //    alpha(1,1)=0;
    //%%%%%%%%%%%%%%%%%%%% alpha forward %%%%%%%%%%%%%%%%%%%%% metric%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%
    //%%%%%%%%%%%%% beta backward metric %%%%%%%%%%%%%% %%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%
    //%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%             
    //             Lezero2=1;
    //       for ii = 1:K
    //           LZ3(1,ii)==2*SNR*x(1,ii)
    //       end
    //       LZ3
    //       asd
    // asd

    for(decoder_fun_fixpt_t_1 = 32'sd0; decoder_fun_fixpt_t_1 <= 32'sd39; decoder_fun_fixpt_t_1 = decoder_fun_fixpt_t_1 + 32'sd1) begin
      decoder_fun_fixpt_LZ[decoder_fun_fixpt_t_1] = 3'sb000;
      decoder_fun_fixpt_Decoded_out[decoder_fun_fixpt_t_1] = 1'b0;
    end


    for(decoder_fun_fixpt_ii_0 = 32'sd0; decoder_fun_fixpt_ii_0 <= 32'sd39; decoder_fun_fixpt_ii_0 = decoder_fun_fixpt_ii_0 + 32'sd1) begin
      decoder_fun_fixpt_add_temp_0[decoder_fun_fixpt_ii_0] = decoder_fun_fixpt_ii_0 + 32'sd1;
      decoder_fun_fixpt_ii = decoder_fun_fixpt_add_temp_0[decoder_fun_fixpt_ii_0][5:0];
      decoder_fun_fixpt_cast[decoder_fun_fixpt_ii_0] = {{3{decoder_fun_fixpt_x[$signed({1'b0, decoder_fun_fixpt_ii}) - 32'sd1][1]}}, {decoder_fun_fixpt_x[$signed({1'b0, decoder_fun_fixpt_ii}) - 32'sd1], 1'b0}};
      decoder_fun_fixpt_LZ[$signed({1'b0, decoder_fun_fixpt_ii}) - 32'sd1] = decoder_fun_fixpt_cast[decoder_fun_fixpt_ii_0][2:0];
      if (decoder_fun_fixpt_LZ[$signed({1'b0, decoder_fun_fixpt_ii}) - 32'sd1] < 3'sb000) begin
        decoder_fun_fixpt_Decoded_out[$signed({1'b0, decoder_fun_fixpt_ii}) - 32'sd1] = 1'b1;
      end
      if (decoder_fun_fixpt_LZ[$signed({1'b0, decoder_fun_fixpt_ii}) - 32'sd1] > 3'sb000) begin
        decoder_fun_fixpt_Decoded_out[$signed({1'b0, decoder_fun_fixpt_ii}) - 32'sd1] = 1'b0;
      end
    end

    //             clc 
    Final_Decoded = decoder_fun_fixpt_Decoded_out;
  end



  assign Final_Decoded_0 = Final_Decoded[0];

  assign Final_Decoded_1 = Final_Decoded[1];

  assign Final_Decoded_2 = Final_Decoded[2];

  assign Final_Decoded_3 = Final_Decoded[3];

  assign Final_Decoded_4 = Final_Decoded[4];

  assign Final_Decoded_5 = Final_Decoded[5];

  assign Final_Decoded_6 = Final_Decoded[6];

  assign Final_Decoded_7 = Final_Decoded[7];

  assign Final_Decoded_8 = Final_Decoded[8];

  assign Final_Decoded_9 = Final_Decoded[9];

  assign Final_Decoded_10 = Final_Decoded[10];

  assign Final_Decoded_11 = Final_Decoded[11];

  assign Final_Decoded_12 = Final_Decoded[12];

  assign Final_Decoded_13 = Final_Decoded[13];

  assign Final_Decoded_14 = Final_Decoded[14];

  assign Final_Decoded_15 = Final_Decoded[15];

  assign Final_Decoded_16 = Final_Decoded[16];

  assign Final_Decoded_17 = Final_Decoded[17];

  assign Final_Decoded_18 = Final_Decoded[18];

  assign Final_Decoded_19 = Final_Decoded[19];

  assign Final_Decoded_20 = Final_Decoded[20];

  assign Final_Decoded_21 = Final_Decoded[21];

  assign Final_Decoded_22 = Final_Decoded[22];

  assign Final_Decoded_23 = Final_Decoded[23];

  assign Final_Decoded_24 = Final_Decoded[24];

  assign Final_Decoded_25 = Final_Decoded[25];

  assign Final_Decoded_26 = Final_Decoded[26];

  assign Final_Decoded_27 = Final_Decoded[27];

  assign Final_Decoded_28 = Final_Decoded[28];

  assign Final_Decoded_29 = Final_Decoded[29];

  assign Final_Decoded_30 = Final_Decoded[30];

  assign Final_Decoded_31 = Final_Decoded[31];

  assign Final_Decoded_32 = Final_Decoded[32];

  assign Final_Decoded_33 = Final_Decoded[33];

  assign Final_Decoded_34 = Final_Decoded[34];

  assign Final_Decoded_35 = Final_Decoded[35];

  assign Final_Decoded_36 = Final_Decoded[36];

  assign Final_Decoded_37 = Final_Decoded[37];

  assign Final_Decoded_38 = Final_Decoded[38];

  assign Final_Decoded_39 = Final_Decoded[39];

endmodule  // decoder_fun_fixpt

